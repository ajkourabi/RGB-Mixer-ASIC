module rgb_led_driver(
    input clk, rst,
    input encoder_A, encoder_B,
    output pwm_red, pwm_green, pwm_blue
);

    
endmodule 